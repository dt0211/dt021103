00168693
00c69693
00168693
01069693
0286a503
00100593
00100613
00158593
00058313
00060393
010000ef
00500633
02c6a623
0140006f
0002f293
007282b3
fff30313
00008067
00000033
